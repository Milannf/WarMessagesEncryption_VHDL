library IEEE;
use IEEE.std_logic_1164.all;

package pattern_pkg is

    subtype PatternStep is std_logic_vector(15 downto 0);
    type PatternArray is array(natural range <>) of PatternStep;

    constant A_PATTERN : PatternArray(0 to 13) := (
        "1111000000000000",
	"1111000000000000",
        "0011110000000000",
	"0011110000000000",
        "0000111100000000",
	"0000111100000000",
        "0000000011110000",
	"0000000011110000",
        "0000000011110000",
	"0000000011110000",
        "0000000000111100",
	"0000000000111100",
        "0000000000011110",
	"0000000000011110"
    );

    constant B_PATTERN : PatternArray(0 to 10) := (
        "1111111111111111",
	"1111111111111111",
        "1110001111000011",
	"1110001111000011",
        "1110001111000011",
	"1110001111000011",
        "1110001111000011",
	"1110001111000011",
        "1111111111111111",
	"1111111111111111",
        "1111111111111111"
    );

    constant C_PATTERN : PatternArray(0 to 8) := (
        "1111111111111111",
	"1111111111111111",
        "1111111111111111",
	"1111000000001111",
        "1111000000001111",
	"1111000000001111",
        "1111000000001111",
	"1111000000001111",
        "1111000000001111"
    );

    constant D_PATTERN : PatternArray(0 to 8) := (
        "1111111111111111",
	"1111111111111111",
        "1110000000000111",
	"1110000000000111",
        "1110000000000111",
	"0011111111111100",
        "0011111111111100",
	"0000111111110000",
        "0000111111110000"
    );

    constant E_PATTERN : PatternArray(0 to 5) := (
        "1111111111111111",
	"1111111111111111",
        "1110000011100011",
	"1110000011100011",
        "1110000011100011",
	"1110000011100011"
    );

    constant F_PATTERN : PatternArray(0 to 5) := (
        "1111111111111111",
	"1111111111111111",
        "0000000011000111",
	"0000000011000111",
        "0000000011000111",
	"0000000011000111"
    );

    constant G_PATTERN : PatternArray(0 to 5) := (
        "1111111111111111",
	"1111111111111111",
        "1111000000001111",
	"1111000000001111",
        "1111000000000000",
	"1111111111100000"
    );

    constant H_PATTERN : PatternArray(0 to 5) := (
        "1111111111111111",
	"1111111111111111",
        "0000000011100000",
	"0000000011100000",
        "1111111111111111",
	"1111111111111111"
    );

    constant I_PATTERN : PatternArray(0 to 2) := (
        "1111111110001111",
	"1111111110001111",
	"1111111110001111"
    );

    constant J_PATTERN : PatternArray(0 to 7) := (
        "1110000000000000",
	"1110000000000000",
        "1110000000000000",
	"1110000000000111",
        "1110000000000111",
	"1110000000000111",
        "1111111111111111",
	"1111111111111111"
    );

    constant K_PATTERN : PatternArray(0 to 5) := (
        "1111111111111111",
	"1111111111111111",
        "0000001111110000",
	"0000001111110000",
        "1111111111001111",
	"1111111111001111"
    );

    constant L_PATTERN : PatternArray(0 to 5) := (
        "1111111111111111",
	"1111111111111111",
        "1111000000000000",
	"1111000000000000",
        "1111000000000000",
	"1111000000000000"
    );

    constant M_PATTERN : PatternArray(0 to 9) := (
        "1111111111110000","1111111111110000",
        "0000000011110000","0000000011110000",
        "1111111111110000","1111111111110000",
        "0000000011110000","0000000011110000",
        "1111111111110000","1111111111110000"
    );

    constant N_PATTERN : PatternArray(0 to 11) := (
        "1111111111111111","1111111111111111",
        "0000000000001111","0000000000011110",
        "0000000000111100","0000000001111000",
        "0000000011110000","0000000111100000",
        "0000001111000000","1111000000000000",
        "1111111111111111","1111111111111111"
    );

    constant O_PATTERN : PatternArray(0 to 10) := (
        "0000111111110000","0011111111111100",
        "0011111111111100","1111111111111111",
        "1100000000000011","1100000000000011",
        "1100000000000011","1111111111111111",
        "0011111111111100","0011111111111100",
        "0000111111110000"
    );

    constant P_PATTERN : PatternArray(0 to 5) := (
        "1111111111111111","1111111111111111",
        "0000000000110001","0000000000110001",
        "0000000000110001","0000000001111111"
    );

    constant Q_PATTERN : PatternArray(0 to 6) := (
        "1111111111111111","1111111111111111",
        "1111100000000011","1001100000000011",
        "1001100000000011","1001111111111111",
        "1001111111111111"
    );

    constant R_PATTERN : PatternArray(0 to 5) := (
        "1111111111111111","1111111111111111",
        "0000000111110011","0000000111110011",
        "1111110011000011","1111110011111111"
    );

    constant S_PATTERN : PatternArray(0 to 5) := (
        "1110001111111111","1110001111111111",
        "1110001110001111","1110001110001111",
        "1111111110001111","1111111110001111"
    );

    constant T_PATTERN : PatternArray(0 to 9) := (
        "0000000000000111","0000000000000111",
        "0000000000000111","0000000000000111",
        "1111111111111111","1111111111111111",
        "0000000000000111","0000000000000111",
        "0000000000000111","0000000000000111"
    );

    constant U_PATTERN : PatternArray(0 to 7) := (
        "1111111111111111","1111111111111111",
        "1110000000000000","1110000000000000",
        "1110000000000000","1110000000000000",
        "1111111111111111","1111111111111111"
    );

    constant V_PATTERN : PatternArray(0 to 12) := (
        "0000000000001111","0000000000001111",
        "0000000011111000","0000000011111000",
        "0011111000000000","0011111000000000",
        "1100000000000000","1100000000000000",
        "0011111000000000","0011111000000000",
        "0000000011111000","0000000011111000",
        "0000000000001111"
    );

    constant W_PATTERN : PatternArray(0 to 9) := (
        "1111111111111100","1111111111111100",
        "1110000000000000","1110000000000000",
        "1111111111111100","1111111111111100",
        "1110000000000000","1110000000000000",
        "1111111111111100","1111111111111100"
    );

    constant X_PATTERN : PatternArray(0 to 9) := (
        "1111000000011111","1111000000011111",
        "0000011100110000","0000011100110000",
        "0000001100000000","0000001100000000",
        "0000011100110000","0000011100110000",
        "1111000000011111","1111000000011111"
    );

    constant Y_PATTERN : PatternArray(0 to 5) := (
        "0000000000111111","0000000000111111",
        "1111111111000000","1111111111000000",
        "0000000000111111","0000000000111111"
    );

    constant Z_PATTERN : PatternArray(0 to 7) := (
        "1110001110000111","1110001110000111",
        "1110001111000111","1110001111000111",
        "1110000001100111","1110000001100111",
        "1110000011000111","1110000011000111"
    );

    constant ZERO_PATTERN : PatternArray(0 to 7) := (
        "0000000000000000","0000000000000000",
        "0000000000000000","0000000000000000",
        "0000000000000000","0000000000000000",
        "0000000000000000","0000000000000000"
    );

end package;

package body pattern_pkg is
end package body;

